// FIFO Package 4
package shared_pkg;           

bit test_finished;  // signal refer to the end of the test bench

// counters declaration
int error_count, correct_count;

endpackage 