package FIFO_shared_pkg;
integer error_count=0;
integer correct_count=0;
    
endpackage